// DE0_Nano_SOPC.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module DE0_Nano_SOPC (
		input  wire        UART_RXD_to_the_RS232_0,                   //                  RS232_0_conduit_end.export
		output wire        UART_TXD_from_the_RS232_0,                 //                RS232_0_conduit_end_1.export
		input  wire        adc_controller_0_conduit_end_sys_clk,      //         adc_controller_0_conduit_end.sys_clk
		output wire        adc_controller_0_conduit_end_ADC_CONVST,   //                                     .ADC_CONVST
		output wire        adc_controller_0_conduit_end_ADC_SDI,      //                                     .ADC_SDI
		output wire        adc_controller_0_conduit_end_ADC_SCK,      //                                     .ADC_SCK
		input  wire        adc_controller_0_conduit_end_ADC_SDO,      //                                     .ADC_SDO
		input  wire        clk_50,                                    //                        clk_50_clk_in.clk
		input  wire        reset_n,                                   //                  clk_50_clk_in_reset.reset_n
		input  wire [1:0]  in_port_to_the_key,                        //              key_external_connection.export
		output wire [7:0]  out_port_from_the_led,                     //              led_external_connection.export
		output wire [31:0] GPIO_out_from_the_motor_controller_0,      //       motor_controller_0_conduit_end.export
		output wire        pll_0_locked_export,                       //                         pll_0_locked.export
		output wire        pll_0_outclk1_clk,                         //                        pll_0_outclk1.clk
		output wire        pll_0_outclk3_clk,                         //                        pll_0_outclk3.clk
		output wire        pll_adc_clk,                               //                              pll_adc.clk
		output wire        pll_io_clk,                                //                               pll_io.clk
		output wire        pll_sys_clk,                               //                              pll_sys.clk
		output wire        kill_sw_from_the_power_management_slave_0, // power_management_slave_0_conduit_end.kill_sw
		output wire [2:0]  mux_from_the_power_management_slave_0,     //                                     .mux
		input  wire        data_to_the_power_management_slave_0,      //                                     .data
		input  wire [3:0]  in_port_to_the_sw                          //               sw_external_connection.export
	);

	wire  [31:0] nios2_gen2_0_data_master_readdata;                                    // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                                 // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                                 // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [24:0] nios2_gen2_0_data_master_address;                                     // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                                  // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                                        // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                                       // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                                   // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                             // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                          // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [24:0] nios2_gen2_0_instruction_master_address;                              // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                                 // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;             // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;               // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;            // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;              // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_motor_controller_0_avalon_slave_0_chipselect;       // mm_interconnect_0:motor_controller_0_avalon_slave_0_chipselect -> motor_controller_0:chipselect
	wire   [4:0] mm_interconnect_0_motor_controller_0_avalon_slave_0_address;          // mm_interconnect_0:motor_controller_0_avalon_slave_0_address -> motor_controller_0:addr
	wire         mm_interconnect_0_motor_controller_0_avalon_slave_0_write;            // mm_interconnect_0:motor_controller_0_avalon_slave_0_write -> motor_controller_0:write
	wire  [31:0] mm_interconnect_0_motor_controller_0_avalon_slave_0_writedata;        // mm_interconnect_0:motor_controller_0_avalon_slave_0_writedata -> motor_controller_0:writedata
	wire         mm_interconnect_0_power_management_slave_0_avalon_slave_0_chipselect; // mm_interconnect_0:power_management_slave_0_avalon_slave_0_chipselect -> power_management_slave_0:chipselect
	wire  [31:0] mm_interconnect_0_power_management_slave_0_avalon_slave_0_readdata;   // power_management_slave_0:readdata -> mm_interconnect_0:power_management_slave_0_avalon_slave_0_readdata
	wire         mm_interconnect_0_power_management_slave_0_avalon_slave_0_read;       // mm_interconnect_0:power_management_slave_0_avalon_slave_0_read -> power_management_slave_0:read
	wire         mm_interconnect_0_power_management_slave_0_avalon_slave_0_write;      // mm_interconnect_0:power_management_slave_0_avalon_slave_0_write -> power_management_slave_0:write
	wire  [31:0] mm_interconnect_0_power_management_slave_0_avalon_slave_0_writedata;  // mm_interconnect_0:power_management_slave_0_avalon_slave_0_writedata -> power_management_slave_0:writedata
	wire         mm_interconnect_0_rs232_0_avalon_slave_0_chipselect;                  // mm_interconnect_0:RS232_0_avalon_slave_0_chipselect -> RS232_0:chipselect
	wire  [31:0] mm_interconnect_0_rs232_0_avalon_slave_0_readdata;                    // RS232_0:readdata -> mm_interconnect_0:RS232_0_avalon_slave_0_readdata
	wire   [0:0] mm_interconnect_0_rs232_0_avalon_slave_0_address;                     // mm_interconnect_0:RS232_0_avalon_slave_0_address -> RS232_0:address
	wire         mm_interconnect_0_rs232_0_avalon_slave_0_read;                        // mm_interconnect_0:RS232_0_avalon_slave_0_read -> RS232_0:read
	wire   [3:0] mm_interconnect_0_rs232_0_avalon_slave_0_byteenable;                  // mm_interconnect_0:RS232_0_avalon_slave_0_byteenable -> RS232_0:byteenable
	wire         mm_interconnect_0_rs232_0_avalon_slave_0_write;                       // mm_interconnect_0:RS232_0_avalon_slave_0_write -> RS232_0:write
	wire  [31:0] mm_interconnect_0_rs232_0_avalon_slave_0_writedata;                   // mm_interconnect_0:RS232_0_avalon_slave_0_writedata -> RS232_0:writedata
	wire         mm_interconnect_0_adc_controller_0_avalon_slave_0_chipselect;         // mm_interconnect_0:adc_controller_0_avalon_slave_0_chipselect -> adc_controller_0:chipselect
	wire  [31:0] mm_interconnect_0_adc_controller_0_avalon_slave_0_readdata;           // adc_controller_0:readdata -> mm_interconnect_0:adc_controller_0_avalon_slave_0_readdata
	wire         mm_interconnect_0_adc_controller_0_avalon_slave_0_read;               // mm_interconnect_0:adc_controller_0_avalon_slave_0_read -> adc_controller_0:read
	wire   [3:0] mm_interconnect_0_adc_controller_0_avalon_slave_0_writebyteenable;    // mm_interconnect_0:adc_controller_0_avalon_slave_0_writebyteenable -> adc_controller_0:addr
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;              // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;           // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;           // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;               // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;                  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;            // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;                 // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;             // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_clock_crossing_io_s0_readdata;                      // clock_crossing_io:s0_readdata -> mm_interconnect_0:clock_crossing_io_s0_readdata
	wire         mm_interconnect_0_clock_crossing_io_s0_waitrequest;                   // clock_crossing_io:s0_waitrequest -> mm_interconnect_0:clock_crossing_io_s0_waitrequest
	wire         mm_interconnect_0_clock_crossing_io_s0_debugaccess;                   // mm_interconnect_0:clock_crossing_io_s0_debugaccess -> clock_crossing_io:s0_debugaccess
	wire   [6:0] mm_interconnect_0_clock_crossing_io_s0_address;                       // mm_interconnect_0:clock_crossing_io_s0_address -> clock_crossing_io:s0_address
	wire         mm_interconnect_0_clock_crossing_io_s0_read;                          // mm_interconnect_0:clock_crossing_io_s0_read -> clock_crossing_io:s0_read
	wire   [3:0] mm_interconnect_0_clock_crossing_io_s0_byteenable;                    // mm_interconnect_0:clock_crossing_io_s0_byteenable -> clock_crossing_io:s0_byteenable
	wire         mm_interconnect_0_clock_crossing_io_s0_readdatavalid;                 // clock_crossing_io:s0_readdatavalid -> mm_interconnect_0:clock_crossing_io_s0_readdatavalid
	wire         mm_interconnect_0_clock_crossing_io_s0_write;                         // mm_interconnect_0:clock_crossing_io_s0_write -> clock_crossing_io:s0_write
	wire  [31:0] mm_interconnect_0_clock_crossing_io_s0_writedata;                     // mm_interconnect_0:clock_crossing_io_s0_writedata -> clock_crossing_io:s0_writedata
	wire   [0:0] mm_interconnect_0_clock_crossing_io_s0_burstcount;                    // mm_interconnect_0:clock_crossing_io_s0_burstcount -> clock_crossing_io:s0_burstcount
	wire         mm_interconnect_0_controller_interrupt_counter_s1_chipselect;         // mm_interconnect_0:controller_interrupt_counter_s1_chipselect -> controller_interrupt_counter:chipselect
	wire  [15:0] mm_interconnect_0_controller_interrupt_counter_s1_readdata;           // controller_interrupt_counter:readdata -> mm_interconnect_0:controller_interrupt_counter_s1_readdata
	wire   [2:0] mm_interconnect_0_controller_interrupt_counter_s1_address;            // mm_interconnect_0:controller_interrupt_counter_s1_address -> controller_interrupt_counter:address
	wire         mm_interconnect_0_controller_interrupt_counter_s1_write;              // mm_interconnect_0:controller_interrupt_counter_s1_write -> controller_interrupt_counter:write_n
	wire  [15:0] mm_interconnect_0_controller_interrupt_counter_s1_writedata;          // mm_interconnect_0:controller_interrupt_counter_s1_writedata -> controller_interrupt_counter:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;                     // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [15:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                       // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [17:0] mm_interconnect_0_onchip_memory2_0_s1_address;                        // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [1:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                     // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                          // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [15:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                      // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                          // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         clock_crossing_io_m0_waitrequest;                                     // mm_interconnect_1:clock_crossing_io_m0_waitrequest -> clock_crossing_io:m0_waitrequest
	wire  [31:0] clock_crossing_io_m0_readdata;                                        // mm_interconnect_1:clock_crossing_io_m0_readdata -> clock_crossing_io:m0_readdata
	wire         clock_crossing_io_m0_debugaccess;                                     // clock_crossing_io:m0_debugaccess -> mm_interconnect_1:clock_crossing_io_m0_debugaccess
	wire   [6:0] clock_crossing_io_m0_address;                                         // clock_crossing_io:m0_address -> mm_interconnect_1:clock_crossing_io_m0_address
	wire         clock_crossing_io_m0_read;                                            // clock_crossing_io:m0_read -> mm_interconnect_1:clock_crossing_io_m0_read
	wire   [3:0] clock_crossing_io_m0_byteenable;                                      // clock_crossing_io:m0_byteenable -> mm_interconnect_1:clock_crossing_io_m0_byteenable
	wire         clock_crossing_io_m0_readdatavalid;                                   // mm_interconnect_1:clock_crossing_io_m0_readdatavalid -> clock_crossing_io:m0_readdatavalid
	wire  [31:0] clock_crossing_io_m0_writedata;                                       // clock_crossing_io:m0_writedata -> mm_interconnect_1:clock_crossing_io_m0_writedata
	wire         clock_crossing_io_m0_write;                                           // clock_crossing_io:m0_write -> mm_interconnect_1:clock_crossing_io_m0_write
	wire   [0:0] clock_crossing_io_m0_burstcount;                                      // clock_crossing_io:m0_burstcount -> mm_interconnect_1:clock_crossing_io_m0_burstcount
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;                       // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;                        // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire         mm_interconnect_1_key_s1_chipselect;                                  // mm_interconnect_1:key_s1_chipselect -> key:chipselect
	wire  [31:0] mm_interconnect_1_key_s1_readdata;                                    // key:readdata -> mm_interconnect_1:key_s1_readdata
	wire   [1:0] mm_interconnect_1_key_s1_address;                                     // mm_interconnect_1:key_s1_address -> key:address
	wire         mm_interconnect_1_key_s1_write;                                       // mm_interconnect_1:key_s1_write -> key:write_n
	wire  [31:0] mm_interconnect_1_key_s1_writedata;                                   // mm_interconnect_1:key_s1_writedata -> key:writedata
	wire         mm_interconnect_1_led_s1_chipselect;                                  // mm_interconnect_1:led_s1_chipselect -> led:chipselect
	wire  [31:0] mm_interconnect_1_led_s1_readdata;                                    // led:readdata -> mm_interconnect_1:led_s1_readdata
	wire   [1:0] mm_interconnect_1_led_s1_address;                                     // mm_interconnect_1:led_s1_address -> led:address
	wire         mm_interconnect_1_led_s1_write;                                       // mm_interconnect_1:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_1_led_s1_writedata;                                   // mm_interconnect_1:led_s1_writedata -> led:writedata
	wire         mm_interconnect_1_sw_s1_chipselect;                                   // mm_interconnect_1:sw_s1_chipselect -> sw:chipselect
	wire  [31:0] mm_interconnect_1_sw_s1_readdata;                                     // sw:readdata -> mm_interconnect_1:sw_s1_readdata
	wire   [1:0] mm_interconnect_1_sw_s1_address;                                      // mm_interconnect_1:sw_s1_address -> sw:address
	wire         mm_interconnect_1_sw_s1_write;                                        // mm_interconnect_1:sw_s1_write -> sw:write_n
	wire  [31:0] mm_interconnect_1_sw_s1_writedata;                                    // mm_interconnect_1:sw_s1_writedata -> sw:writedata
	wire         irq_mapper_receiver3_irq;                                             // jtag_uart:av_irq -> irq_mapper:receiver3_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                                 // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         irq_mapper_receiver0_irq;                                             // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                        // power_management_slave_0:error -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver1_irq;                                             // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                                    // RS232_0:irq -> irq_synchronizer_001:receiver_irq
	wire         irq_mapper_receiver2_irq;                                             // irq_synchronizer_002:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_002_receiver_irq;                                    // controller_interrupt_counter:irq -> irq_synchronizer_002:receiver_irq
	wire         irq_mapper_receiver4_irq;                                             // irq_synchronizer_003:sender_irq -> irq_mapper:receiver4_irq
	wire   [0:0] irq_synchronizer_003_receiver_irq;                                    // key:irq -> irq_synchronizer_003:receiver_irq
	wire         irq_mapper_receiver5_irq;                                             // irq_synchronizer_004:sender_irq -> irq_mapper:receiver5_irq
	wire   [0:0] irq_synchronizer_004_receiver_irq;                                    // sw:irq -> irq_synchronizer_004:receiver_irq
	wire         rst_controller_reset_out_reset;                                       // rst_controller:reset_out -> [RS232_0:reset, controller_interrupt_counter:reset_n, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, mm_interconnect_0:motor_controller_0_reset_reset_bridge_in_reset_reset, motor_controller_0:reset, power_management_slave_0:reset]
	wire         nios2_gen2_0_debug_reset_request_reset;                               // nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1, rst_controller_003:reset_in1]
	wire         rst_controller_001_reset_out_reset;                                   // rst_controller_001:reset_out -> [adc_controller_0:spi_reset, mm_interconnect_0:adc_controller_0_reset_sink_reset_bridge_in_reset_reset]
	wire         rst_controller_002_reset_out_reset;                                   // rst_controller_002:reset_out -> [clock_crossing_io:m0_reset, irq_synchronizer_003:receiver_reset, irq_synchronizer_004:receiver_reset, key:reset_n, led:reset_n, mm_interconnect_1:clock_crossing_io_m0_reset_reset_bridge_in_reset_reset, sw:reset_n, sysid:reset_n]
	wire         rst_controller_003_reset_out_reset;                                   // rst_controller_003:reset_out -> [clock_crossing_io:s0_reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, irq_synchronizer_004:sender_reset, jtag_uart:rst_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_memory2_0:reset, rst_translator:in_reset]
	wire         rst_controller_003_reset_out_reset_req;                               // rst_controller_003:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]

	Altera_UP_Avalon_RS232 rs232_0 (
		.clk        (clk_50),                                              //            clock.clk
		.reset      (rst_controller_reset_out_reset),                      //            reset.reset
		.address    (mm_interconnect_0_rs232_0_avalon_slave_0_address),    //   avalon_slave_0.address
		.chipselect (mm_interconnect_0_rs232_0_avalon_slave_0_chipselect), //                 .chipselect
		.byteenable (mm_interconnect_0_rs232_0_avalon_slave_0_byteenable), //                 .byteenable
		.read       (mm_interconnect_0_rs232_0_avalon_slave_0_read),       //                 .read
		.write      (mm_interconnect_0_rs232_0_avalon_slave_0_write),      //                 .write
		.writedata  (mm_interconnect_0_rs232_0_avalon_slave_0_writedata),  //                 .writedata
		.readdata   (mm_interconnect_0_rs232_0_avalon_slave_0_readdata),   //                 .readdata
		.UART_RXD   (UART_RXD_to_the_RS232_0),                             //      conduit_end.export
		.UART_TXD   (UART_TXD_from_the_RS232_0),                           //    conduit_end_1.export
		.irq        (irq_synchronizer_001_receiver_irq)                    // interrupt_sender.irq
	);

	adc_controller adc_controller_0 (
		.chipselect (mm_interconnect_0_adc_controller_0_avalon_slave_0_chipselect),       // avalon_slave_0.chipselect
		.addr       (~mm_interconnect_0_adc_controller_0_avalon_slave_0_writebyteenable), //               .writebyteenable_n
		.read       (mm_interconnect_0_adc_controller_0_avalon_slave_0_read),             //               .read
		.readdata   (mm_interconnect_0_adc_controller_0_avalon_slave_0_readdata),         //               .readdata
		.sys_clk    (adc_controller_0_conduit_end_sys_clk),                               //    conduit_end.export
		.ADC_CONVST (adc_controller_0_conduit_end_ADC_CONVST),                            //               .export
		.ADC_SDI    (adc_controller_0_conduit_end_ADC_SDI),                               //               .export
		.ADC_SCK    (adc_controller_0_conduit_end_ADC_SCK),                               //               .export
		.ADC_SDO    (adc_controller_0_conduit_end_ADC_SDO),                               //               .export
		.spi_clk    (pll_adc_clk),                                                        //     clock_sink.clk
		.spi_reset  (rst_controller_001_reset_out_reset)                                  //     reset_sink.reset
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (7),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (16),
		.RESPONSE_FIFO_DEPTH (32),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) clock_crossing_io (
		.m0_clk           (pll_io_clk),                                           //   m0_clk.clk
		.m0_reset         (rst_controller_002_reset_out_reset),                   // m0_reset.reset
		.s0_clk           (pll_sys_clk),                                          //   s0_clk.clk
		.s0_reset         (rst_controller_003_reset_out_reset),                   // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_clock_crossing_io_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_clock_crossing_io_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_clock_crossing_io_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_clock_crossing_io_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_clock_crossing_io_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_clock_crossing_io_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_clock_crossing_io_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_clock_crossing_io_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_clock_crossing_io_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_clock_crossing_io_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (clock_crossing_io_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (clock_crossing_io_m0_readdata),                        //         .readdata
		.m0_readdatavalid (clock_crossing_io_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (clock_crossing_io_m0_burstcount),                      //         .burstcount
		.m0_writedata     (clock_crossing_io_m0_writedata),                       //         .writedata
		.m0_address       (clock_crossing_io_m0_address),                         //         .address
		.m0_write         (clock_crossing_io_m0_write),                           //         .write
		.m0_read          (clock_crossing_io_m0_read),                            //         .read
		.m0_byteenable    (clock_crossing_io_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (clock_crossing_io_m0_debugaccess)                      //         .debugaccess
	);

	DE0_Nano_SOPC_controller_interrupt_counter controller_interrupt_counter (
		.clk        (clk_50),                                                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                              // reset.reset_n
		.address    (mm_interconnect_0_controller_interrupt_counter_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_controller_interrupt_counter_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_controller_interrupt_counter_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_controller_interrupt_counter_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_controller_interrupt_counter_s1_write),     //      .write_n
		.irq        (irq_synchronizer_002_receiver_irq)                             //   irq.irq
	);

	DE0_Nano_SOPC_jtag_uart jtag_uart (
		.clk            (pll_sys_clk),                                               //               clk.clk
		.rst_n          (~rst_controller_003_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver3_irq)                                   //               irq.irq
	);

	DE0_Nano_SOPC_key key (
		.clk        (pll_io_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_1_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_key_s1_readdata),   //                    .readdata
		.in_port    (in_port_to_the_key),                  // external_connection.export
		.irq        (irq_synchronizer_003_receiver_irq)    //                 irq.irq
	);

	DE0_Nano_SOPC_led led (
		.clk        (pll_io_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_1_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_s1_readdata),   //                    .readdata
		.out_port   (out_port_from_the_led)                // external_connection.export
	);

	slave_controller motor_controller_0 (
		.clk        (clk_50),                                                         //          clock.clk
		.chipselect (mm_interconnect_0_motor_controller_0_avalon_slave_0_chipselect), // avalon_slave_0.chipselect
		.write      (mm_interconnect_0_motor_controller_0_avalon_slave_0_write),      //               .write
		.addr       (mm_interconnect_0_motor_controller_0_avalon_slave_0_address),    //               .address
		.writedata  (mm_interconnect_0_motor_controller_0_avalon_slave_0_writedata),  //               .writedata
		.GPIO_out   (GPIO_out_from_the_motor_controller_0),                           //    conduit_end.export
		.reset      (rst_controller_reset_out_reset)                                  //          reset.reset
	);

	DE0_Nano_SOPC_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (pll_sys_clk),                                                //                       clk.clk
		.reset_n                             (~rst_controller_003_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_003_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	DE0_Nano_SOPC_onchip_memory2_0 onchip_memory2_0 (
		.clk        (pll_sys_clk),                                      //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_003_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_003_reset_out_reset_req)            //       .reset_req
	);

	DE0_Nano_SOPC_pll_0 pll_0 (
		.refclk   (clk_50),              //  refclk.clk
		.rst      (~reset_n),            //   reset.reset
		.outclk_0 (pll_sys_clk),         // outclk0.clk
		.outclk_1 (pll_0_outclk1_clk),   // outclk1.clk
		.outclk_2 (pll_io_clk),          // outclk2.clk
		.outclk_3 (pll_0_outclk3_clk),   // outclk3.clk
		.outclk_4 (pll_adc_clk),         // outclk4.clk
		.locked   (pll_0_locked_export)  //  locked.export
	);

	power_management_slave power_management_slave_0 (
		.chipselect (mm_interconnect_0_power_management_slave_0_avalon_slave_0_chipselect), //   avalon_slave_0.chipselect
		.write      (mm_interconnect_0_power_management_slave_0_avalon_slave_0_write),      //                 .write
		.read       (mm_interconnect_0_power_management_slave_0_avalon_slave_0_read),       //                 .read
		.writedata  (mm_interconnect_0_power_management_slave_0_avalon_slave_0_writedata),  //                 .writedata
		.readdata   (mm_interconnect_0_power_management_slave_0_avalon_slave_0_readdata),   //                 .readdata
		.clk        (clk_50),                                                               //            clock.clk
		.kill_sw    (kill_sw_from_the_power_management_slave_0),                            //      conduit_end.export
		.mux        (mux_from_the_power_management_slave_0),                                //                 .export
		.data       (data_to_the_power_management_slave_0),                                 //                 .export
		.error      (irq_synchronizer_receiver_irq),                                        // interrupt_sender.irq
		.reset      (rst_controller_reset_out_reset)                                        //            reset.reset
	);

	DE0_Nano_SOPC_sw sw (
		.clk        (pll_io_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_1_sw_s1_address),     //                  s1.address
		.write_n    (~mm_interconnect_1_sw_s1_write),      //                    .write_n
		.writedata  (mm_interconnect_1_sw_s1_writedata),   //                    .writedata
		.chipselect (mm_interconnect_1_sw_s1_chipselect),  //                    .chipselect
		.readdata   (mm_interconnect_1_sw_s1_readdata),    //                    .readdata
		.in_port    (in_port_to_the_sw),                   // external_connection.export
		.irq        (irq_synchronizer_004_receiver_irq)    //                 irq.irq
	);

	DE0_Nano_SOPC_sysid sysid (
		.clock    (pll_io_clk),                                     //           clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	DE0_Nano_SOPC_mm_interconnect_0 mm_interconnect_0 (
		.clk_50_clk_clk                                          (clk_50),                                                               //                                        clk_50_clk.clk
		.pll_0_outclk0_clk                                       (pll_sys_clk),                                                          //                                     pll_0_outclk0.clk
		.pll_0_outclk4_clk                                       (pll_adc_clk),                                                          //                                     pll_0_outclk4.clk
		.adc_controller_0_reset_sink_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                                   // adc_controller_0_reset_sink_reset_bridge_in_reset.reset
		.motor_controller_0_reset_reset_bridge_in_reset_reset    (rst_controller_reset_out_reset),                                       //    motor_controller_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset          (rst_controller_003_reset_out_reset),                                   //          nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address                        (nios2_gen2_0_data_master_address),                                     //                          nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                    (nios2_gen2_0_data_master_waitrequest),                                 //                                                  .waitrequest
		.nios2_gen2_0_data_master_byteenable                     (nios2_gen2_0_data_master_byteenable),                                  //                                                  .byteenable
		.nios2_gen2_0_data_master_read                           (nios2_gen2_0_data_master_read),                                        //                                                  .read
		.nios2_gen2_0_data_master_readdata                       (nios2_gen2_0_data_master_readdata),                                    //                                                  .readdata
		.nios2_gen2_0_data_master_write                          (nios2_gen2_0_data_master_write),                                       //                                                  .write
		.nios2_gen2_0_data_master_writedata                      (nios2_gen2_0_data_master_writedata),                                   //                                                  .writedata
		.nios2_gen2_0_data_master_debugaccess                    (nios2_gen2_0_data_master_debugaccess),                                 //                                                  .debugaccess
		.nios2_gen2_0_instruction_master_address                 (nios2_gen2_0_instruction_master_address),                              //                   nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest             (nios2_gen2_0_instruction_master_waitrequest),                          //                                                  .waitrequest
		.nios2_gen2_0_instruction_master_read                    (nios2_gen2_0_instruction_master_read),                                 //                                                  .read
		.nios2_gen2_0_instruction_master_readdata                (nios2_gen2_0_instruction_master_readdata),                             //                                                  .readdata
		.adc_controller_0_avalon_slave_0_read                    (mm_interconnect_0_adc_controller_0_avalon_slave_0_read),               //                   adc_controller_0_avalon_slave_0.read
		.adc_controller_0_avalon_slave_0_readdata                (mm_interconnect_0_adc_controller_0_avalon_slave_0_readdata),           //                                                  .readdata
		.adc_controller_0_avalon_slave_0_writebyteenable         (mm_interconnect_0_adc_controller_0_avalon_slave_0_writebyteenable),    //                                                  .writebyteenable
		.adc_controller_0_avalon_slave_0_chipselect              (mm_interconnect_0_adc_controller_0_avalon_slave_0_chipselect),         //                                                  .chipselect
		.clock_crossing_io_s0_address                            (mm_interconnect_0_clock_crossing_io_s0_address),                       //                              clock_crossing_io_s0.address
		.clock_crossing_io_s0_write                              (mm_interconnect_0_clock_crossing_io_s0_write),                         //                                                  .write
		.clock_crossing_io_s0_read                               (mm_interconnect_0_clock_crossing_io_s0_read),                          //                                                  .read
		.clock_crossing_io_s0_readdata                           (mm_interconnect_0_clock_crossing_io_s0_readdata),                      //                                                  .readdata
		.clock_crossing_io_s0_writedata                          (mm_interconnect_0_clock_crossing_io_s0_writedata),                     //                                                  .writedata
		.clock_crossing_io_s0_burstcount                         (mm_interconnect_0_clock_crossing_io_s0_burstcount),                    //                                                  .burstcount
		.clock_crossing_io_s0_byteenable                         (mm_interconnect_0_clock_crossing_io_s0_byteenable),                    //                                                  .byteenable
		.clock_crossing_io_s0_readdatavalid                      (mm_interconnect_0_clock_crossing_io_s0_readdatavalid),                 //                                                  .readdatavalid
		.clock_crossing_io_s0_waitrequest                        (mm_interconnect_0_clock_crossing_io_s0_waitrequest),                   //                                                  .waitrequest
		.clock_crossing_io_s0_debugaccess                        (mm_interconnect_0_clock_crossing_io_s0_debugaccess),                   //                                                  .debugaccess
		.controller_interrupt_counter_s1_address                 (mm_interconnect_0_controller_interrupt_counter_s1_address),            //                   controller_interrupt_counter_s1.address
		.controller_interrupt_counter_s1_write                   (mm_interconnect_0_controller_interrupt_counter_s1_write),              //                                                  .write
		.controller_interrupt_counter_s1_readdata                (mm_interconnect_0_controller_interrupt_counter_s1_readdata),           //                                                  .readdata
		.controller_interrupt_counter_s1_writedata               (mm_interconnect_0_controller_interrupt_counter_s1_writedata),          //                                                  .writedata
		.controller_interrupt_counter_s1_chipselect              (mm_interconnect_0_controller_interrupt_counter_s1_chipselect),         //                                                  .chipselect
		.jtag_uart_avalon_jtag_slave_address                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),                //                       jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                  //                                                  .write
		.jtag_uart_avalon_jtag_slave_read                        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                   //                                                  .read
		.jtag_uart_avalon_jtag_slave_readdata                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),               //                                                  .readdata
		.jtag_uart_avalon_jtag_slave_writedata                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),              //                                                  .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),            //                                                  .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),             //                                                  .chipselect
		.motor_controller_0_avalon_slave_0_address               (mm_interconnect_0_motor_controller_0_avalon_slave_0_address),          //                 motor_controller_0_avalon_slave_0.address
		.motor_controller_0_avalon_slave_0_write                 (mm_interconnect_0_motor_controller_0_avalon_slave_0_write),            //                                                  .write
		.motor_controller_0_avalon_slave_0_writedata             (mm_interconnect_0_motor_controller_0_avalon_slave_0_writedata),        //                                                  .writedata
		.motor_controller_0_avalon_slave_0_chipselect            (mm_interconnect_0_motor_controller_0_avalon_slave_0_chipselect),       //                                                  .chipselect
		.nios2_gen2_0_debug_mem_slave_address                    (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),               //                      nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                      (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),                 //                                                  .write
		.nios2_gen2_0_debug_mem_slave_read                       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),                  //                                                  .read
		.nios2_gen2_0_debug_mem_slave_readdata                   (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),              //                                                  .readdata
		.nios2_gen2_0_debug_mem_slave_writedata                  (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),             //                                                  .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable                 (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),            //                                                  .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),           //                                                  .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),           //                                                  .debugaccess
		.onchip_memory2_0_s1_address                             (mm_interconnect_0_onchip_memory2_0_s1_address),                        //                               onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                               (mm_interconnect_0_onchip_memory2_0_s1_write),                          //                                                  .write
		.onchip_memory2_0_s1_readdata                            (mm_interconnect_0_onchip_memory2_0_s1_readdata),                       //                                                  .readdata
		.onchip_memory2_0_s1_writedata                           (mm_interconnect_0_onchip_memory2_0_s1_writedata),                      //                                                  .writedata
		.onchip_memory2_0_s1_byteenable                          (mm_interconnect_0_onchip_memory2_0_s1_byteenable),                     //                                                  .byteenable
		.onchip_memory2_0_s1_chipselect                          (mm_interconnect_0_onchip_memory2_0_s1_chipselect),                     //                                                  .chipselect
		.onchip_memory2_0_s1_clken                               (mm_interconnect_0_onchip_memory2_0_s1_clken),                          //                                                  .clken
		.power_management_slave_0_avalon_slave_0_write           (mm_interconnect_0_power_management_slave_0_avalon_slave_0_write),      //           power_management_slave_0_avalon_slave_0.write
		.power_management_slave_0_avalon_slave_0_read            (mm_interconnect_0_power_management_slave_0_avalon_slave_0_read),       //                                                  .read
		.power_management_slave_0_avalon_slave_0_readdata        (mm_interconnect_0_power_management_slave_0_avalon_slave_0_readdata),   //                                                  .readdata
		.power_management_slave_0_avalon_slave_0_writedata       (mm_interconnect_0_power_management_slave_0_avalon_slave_0_writedata),  //                                                  .writedata
		.power_management_slave_0_avalon_slave_0_chipselect      (mm_interconnect_0_power_management_slave_0_avalon_slave_0_chipselect), //                                                  .chipselect
		.RS232_0_avalon_slave_0_address                          (mm_interconnect_0_rs232_0_avalon_slave_0_address),                     //                            RS232_0_avalon_slave_0.address
		.RS232_0_avalon_slave_0_write                            (mm_interconnect_0_rs232_0_avalon_slave_0_write),                       //                                                  .write
		.RS232_0_avalon_slave_0_read                             (mm_interconnect_0_rs232_0_avalon_slave_0_read),                        //                                                  .read
		.RS232_0_avalon_slave_0_readdata                         (mm_interconnect_0_rs232_0_avalon_slave_0_readdata),                    //                                                  .readdata
		.RS232_0_avalon_slave_0_writedata                        (mm_interconnect_0_rs232_0_avalon_slave_0_writedata),                   //                                                  .writedata
		.RS232_0_avalon_slave_0_byteenable                       (mm_interconnect_0_rs232_0_avalon_slave_0_byteenable),                  //                                                  .byteenable
		.RS232_0_avalon_slave_0_chipselect                       (mm_interconnect_0_rs232_0_avalon_slave_0_chipselect)                   //                                                  .chipselect
	);

	DE0_Nano_SOPC_mm_interconnect_1 mm_interconnect_1 (
		.pll_0_outclk2_clk                                      (pll_io_clk),                                     //                                    pll_0_outclk2.clk
		.clock_crossing_io_m0_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),             // clock_crossing_io_m0_reset_reset_bridge_in_reset.reset
		.clock_crossing_io_m0_address                           (clock_crossing_io_m0_address),                   //                             clock_crossing_io_m0.address
		.clock_crossing_io_m0_waitrequest                       (clock_crossing_io_m0_waitrequest),               //                                                 .waitrequest
		.clock_crossing_io_m0_burstcount                        (clock_crossing_io_m0_burstcount),                //                                                 .burstcount
		.clock_crossing_io_m0_byteenable                        (clock_crossing_io_m0_byteenable),                //                                                 .byteenable
		.clock_crossing_io_m0_read                              (clock_crossing_io_m0_read),                      //                                                 .read
		.clock_crossing_io_m0_readdata                          (clock_crossing_io_m0_readdata),                  //                                                 .readdata
		.clock_crossing_io_m0_readdatavalid                     (clock_crossing_io_m0_readdatavalid),             //                                                 .readdatavalid
		.clock_crossing_io_m0_write                             (clock_crossing_io_m0_write),                     //                                                 .write
		.clock_crossing_io_m0_writedata                         (clock_crossing_io_m0_writedata),                 //                                                 .writedata
		.clock_crossing_io_m0_debugaccess                       (clock_crossing_io_m0_debugaccess),               //                                                 .debugaccess
		.key_s1_address                                         (mm_interconnect_1_key_s1_address),               //                                           key_s1.address
		.key_s1_write                                           (mm_interconnect_1_key_s1_write),                 //                                                 .write
		.key_s1_readdata                                        (mm_interconnect_1_key_s1_readdata),              //                                                 .readdata
		.key_s1_writedata                                       (mm_interconnect_1_key_s1_writedata),             //                                                 .writedata
		.key_s1_chipselect                                      (mm_interconnect_1_key_s1_chipselect),            //                                                 .chipselect
		.led_s1_address                                         (mm_interconnect_1_led_s1_address),               //                                           led_s1.address
		.led_s1_write                                           (mm_interconnect_1_led_s1_write),                 //                                                 .write
		.led_s1_readdata                                        (mm_interconnect_1_led_s1_readdata),              //                                                 .readdata
		.led_s1_writedata                                       (mm_interconnect_1_led_s1_writedata),             //                                                 .writedata
		.led_s1_chipselect                                      (mm_interconnect_1_led_s1_chipselect),            //                                                 .chipselect
		.sw_s1_address                                          (mm_interconnect_1_sw_s1_address),                //                                            sw_s1.address
		.sw_s1_write                                            (mm_interconnect_1_sw_s1_write),                  //                                                 .write
		.sw_s1_readdata                                         (mm_interconnect_1_sw_s1_readdata),               //                                                 .readdata
		.sw_s1_writedata                                        (mm_interconnect_1_sw_s1_writedata),              //                                                 .writedata
		.sw_s1_chipselect                                       (mm_interconnect_1_sw_s1_chipselect),             //                                                 .chipselect
		.sysid_control_slave_address                            (mm_interconnect_1_sysid_control_slave_address),  //                              sysid_control_slave.address
		.sysid_control_slave_readdata                           (mm_interconnect_1_sysid_control_slave_readdata)  //                                                 .readdata
	);

	DE0_Nano_SOPC_irq_mapper irq_mapper (
		.clk           (pll_sys_clk),                        //       clk.clk
		.reset         (rst_controller_003_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),           // receiver5.irq
		.sender_irq    (nios2_gen2_0_irq_irq)                //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clk_50),                             //       receiver_clk.clk
		.sender_clk     (pll_sys_clk),                        //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_003_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (clk_50),                             //       receiver_clk.clk
		.sender_clk     (pll_sys_clk),                        //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_003_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (clk_50),                             //       receiver_clk.clk
		.sender_clk     (pll_sys_clk),                        //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_003_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_003 (
		.receiver_clk   (pll_io_clk),                         //       receiver_clk.clk
		.sender_clk     (pll_sys_clk),                        //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_003_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_003_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver4_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_004 (
		.receiver_clk   (pll_io_clk),                         //       receiver_clk.clk
		.sender_clk     (pll_sys_clk),                        //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_003_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_004_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver5_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_n),                               // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_50),                                 //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_n),                               // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (pll_adc_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_n),                               // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (pll_io_clk),                             //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_n),                               // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (pll_sys_clk),                            //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_003_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
